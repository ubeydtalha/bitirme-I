.PARAM
+ LM1 = 8.936375908806574e-06
+ LM2 = 3.01857225250581e-06
+ LM3 = 9.434686135561626e-06
+ WM1 = 5.273435246069726e-05
+ WM2 = 7.609232643652538e-05
+ WM3 = 8.366153923717727e-05
+ Rb = 22530.274371633714
+ Vb = 0.996996294312359
