.PARAM
+ LM1 = True
+ LM2 = True
+ LM3 = False
+ WM1 = True
+ WM2 = True
+ WM3 = False
+ Rb = False
+ Vb = True
