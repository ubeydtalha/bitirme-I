.PARAM
+ LM1 = True
+ LM2 = True
+ LM3 = True
+ WM1 = False
+ WM2 = True
+ WM3 = True
+ Rb = True
+ Vb = False
