.PARAM
+ LM1 = 8.384567841222737e-06
+ LM2 = 4.272405486964919e-06
+ LM3 = 5.066472271942056e-06
+ WM1 = 2.4944455932182386e-05
+ WM2 = 7.518661159751893e-05
+ WM3 = 5.9928397724459784e-05
+ Rb = 18395.845272340088
+ Vb = 0.4154274159384351
