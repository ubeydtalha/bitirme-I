.PARAM
+ LM1 = 1.0092e-06
+ LM2 = 1.4842e-06
+ LM3 = 1.5565e-06
+ WM1 = 2.1734e-05
+ WM2 = 4.6268e-05
+ WM3 = 6.2646e-05
+ Rb = 10000
+ Vb = 0.55
