.PARAM
+ LM1 = 2.4706530569702892e-06
+ LM2 = 1.9544413255161715e-06
+ LM3 = 6.69255583353073e-07
+ WM1 = 6.0401761205027166e-05
+ WM2 = 4.008350842017432e-05
+ WM3 = 0.00016670954335992028
+ Rb = 18180.468000978275
+ Vb = 0.6842750783987592
